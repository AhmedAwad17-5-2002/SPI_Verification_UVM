interface SPI_if(clk);
	input clk;
	logic MOSI, SS_n,rst_n,MISO,MISO_G;
endinterface : SPI_if